 library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity debouncer is
    port(   clock : in std_logic;
            n_reset : in std_logic;
            button_in : in std_logic;
            pulse_out : out std_logic
        );
end debouncer;

architecture behav of debouncer is

--the below constants decide the working parameters.
--the higher this is, the more longer time the user has to press the button.
constant COUNT_MAX : integer := 100; 
--set it '1' if the button creates a high pulse when its pressed, otherwise '0'.
signal latched_state : std_logic := '1';

signal count : integer := 0;
type state_type is (idle,wait_time); --state machine
signal state : state_type := idle;

begin
  
process(n_reset,clock)
begin
	if(n_reset = '0') then
		
		state <= idle;
		pulse_out <= '0';
	
	elsif(rising_edge(clock)) then
       
		case (state) is
			when idle =>
                
				if(button_in = latched_state) then  
						
					state <= idle; --wait until button is pressed.
				else
					state <= wait_time;

				end if;
			
			when wait_time =>
				 
				if(count = COUNT_MAX) then
					
					count <= 0;
					state <= idle; 
					
					if(button_in /= latched_state) then
						pulse_out <= button_in;
						latched_state <= button_in;
					end if; 
                
				else
					count <= count + 1;
				end if; 
					
			end case;       
    end if;        
end process;                  
                                                                                
end architecture behav;