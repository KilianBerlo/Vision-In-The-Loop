
module first_nios2_system (
	clk_clk,
	reset_reset_n,
	esl_bus_demo_0_user_interface_export);	

	input		clk_clk;
	input		reset_reset_n;
	output	[7:0]	esl_bus_demo_0_user_interface_export;
endmodule
